`define FPGA_MODE 1
