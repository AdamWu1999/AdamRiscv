`timescale 1ns/1ps


module tbtop();

`include "../../testbench/instance"
`include "../../testbench/environment.sv"
`include "../../testbench/ext_behavior_task/simple_task/simple.v"
`include "user.sv"



endmodule
